//#############################################################################
// WRITTEN BY ANNIE (WEI) DAI PLOTTING PRETTY LITTLE PICTURES OF
// A BOX HUMAN MODEL. THIS MODULE RETURNS THE BEGINNING AND ENDING 
// COORDINATES OF A LINE WHICH ARE NEEDED FOR THE BRESENHAM LINE DRAWING MODULE
// SPRING 2013
//#############################################################################
/////////////////////////////////////////////////////
//// UPPER BODY MODEL COORDINATES LOOKUP TABLE///////
/////////////////////////////////////////////////////
module body_LUT(x1,y1,x2,y2,oldhcx,oldhcy,oldlcx,oldlcy,oldrcx,oldrcy,lineCount);
output reg [9:0] x1,x2;
output reg [8:0] y1,y2;
input [5:0] lineCount;
input [9:0] oldhcx,oldhcy,oldlcx,oldlcy,oldrcx,oldrcy;

always @(lineCount)
begin
	case (lineCount)
					6'd0:
					begin
						x1<=(oldhcx)-10'd50;
						y1<=(oldhcy)-9'd10;
						x2<=(oldhcx)+10'd50;
						y2<=(oldhcy)-9'd10;
					end
					6'd1:
					begin
						x1<=(oldhcx)+10'd50;
						y1<=(oldhcy)-9'd10;
						x2<=(oldhcx)+10'd50;
						y2<=(oldhcy)+9'd90;
					end
					6'd2:
					begin
						x1<=(oldhcx)+10'd50;
						y1<=(oldhcy)+9'd90;
						x2<=(oldhcx)-10'd50;
						y2<=(oldhcy)+9'd90;
					end
					6'd3:
					begin
						x1<=(oldhcx)-10'd50;
						y1<=(oldhcy)+9'd90;
						x2<=(oldhcx)-10'd50;
						y2<=(oldhcy)-9'd10;
					end
					6'd4:
					begin
						x1<=(oldhcx)-10'd30+oldhcx[9:3]-6'd40;
						y1<=(oldhcy)+9'd10+oldhcy[8:3]-5'd10;
						x2<=(oldhcx)+10'd30+oldhcx[9:3]-6'd40;
						y2<=(oldhcy)+9'd10+oldhcy[8:3]-5'd10;
					end
					6'd5:
					begin
						x1<=(oldhcx)+10'd30+oldhcx[9:3]-6'd40;
						y1<=(oldhcy)+9'd10+oldhcy[8:3]-5'd10;
						x2<=(oldhcx)+10'd30+oldhcx[9:3]-6'd40;
						y2<=(oldhcy)+9'd70+oldhcy[8:3]-5'd10;
					end
					6'd6:
					begin
						x1<=(oldhcx)+10'd30+oldhcx[9:3]-6'd40;
						y1<=(oldhcy)+9'd70+oldhcy[8:3]-5'd10;
						x2<=(oldhcx)-10'd30+oldhcx[9:3]-6'd40;
						y2<=(oldhcy)+9'd70+oldhcy[8:3]-5'd10;
					end
					6'd7:
					begin
						x1<=(oldhcx)-10'd30+oldhcx[9:3]-6'd40;
						y1<=(oldhcy)+9'd70+oldhcy[8:3]-5'd10;
						x2<=(oldhcx)-10'd30+oldhcx[9:3]-6'd40;
						y2<=(oldhcy)+9'd10+oldhcy[8:3]-5'd10;
					end
					6'd8:
					begin
						x1<=(oldhcx)-10'd30+oldhcx[9:3]-6'd40;
						y1<=(oldhcy)+9'd10+oldhcy[8:3]-5'd10;
						x2<=(oldhcx)-10'd50;
						y2<=(oldhcy)-9'd10;
					end
					6'd9:
					begin
						x1<=(oldhcx)+10'd30+oldhcx[9:3]-6'd40;
						y1<=(oldhcy)+9'd10+oldhcy[8:3]-5'd10;
						x2<=(oldhcx)+10'd50;
						y2<=(oldhcy)-9'd10;
					end
					6'd10:
					begin
						x1<=(oldhcx)+10'd30+oldhcx[9:3]-6'd40;
						y1<=(oldhcy)+9'd70+oldhcy[8:3]-5'd10;
						x2<=(oldhcx)+10'd50;
						y2<=(oldhcy)+9'd90;
					end
					6'd11:
					begin
						x1<=(oldhcx)-10'd30+oldhcx[9:3]-6'd40;
						y1<=(oldhcy)+9'd70+oldhcy[8:3]-5'd10;
						x2<=(oldhcx)-10'd50;
						y2<=(oldhcy)+9'd90;
					end
					6'd12:
					begin
						x1<=oldhcx-10'd80;//horizontal arm top
						y1<=oldhcy+9'd110;
						x2<=oldhcx-10'd60;
						y2<=oldhcy+9'd110;
					end
					6'd13:
					begin
						x1<=oldhcx-10'd80;//armleft
						y1<=oldhcy+9'd110;
						x2<=oldlcx-10'd20;
						y2<=oldlcy;
					end
					6'd14:
					begin
						x1<=oldhcx-10'd60;
						y1<=oldhcy+9'd110;
						x2<=oldlcx+10'd20;
						y2<=oldlcy;
					end
					6'd15:
					begin
						x1<=oldlcx-10'd20;
						y1<=oldlcy;
						x2<=oldlcx+10'd20;
						y2<=oldlcy;
					end
					6'd16:
					begin
						x1<=oldlcx-10'd20;
						y1<=oldlcy;
						x2<=oldlcx-10'd20;
						y2<=oldlcy-oldlcy[8:3]+10'd60;
					end
					6'd17:
					begin
						x1<=oldlcx+10'd20;
						y1<=oldlcy;
						x2<=oldlcx+10'd20;
						y2<=oldlcy-oldlcy[8:3]+10'd60;
					end
					6'd18:
					begin
						x1<=oldlcx-10'd20;
						y1<=oldlcy-oldlcy[8:3]+10'd60;
						x2<=oldlcx+10'd20;
						y2<=oldlcy-oldlcy[8:3]+10'd60;
					end
					6'd19:
					begin
						x1<=oldhcx-10'd80;//horizontal arm top bot
						y1<=oldhcy+9'd130;
						x2<=oldhcx-10'd60;
						y2<=oldhcy+9'd130;
					end
					6'd20:
					begin
						x1<=oldhcx-10'd80;//horizontal arm top bot
						y1<=oldhcy+9'd130;
						x2<=oldlcx-10'd20;
						y2<=oldlcy-oldlcy[8:3]+10'd60;					
					end
					6'd21:
					begin
						x1<=oldhcx-10'd60;
						y1<=oldhcy+9'd130;
						x2<=oldlcx+10'd20;
						y2<=oldlcy-oldlcy[8:3]+10'd60;
					end
					6'd22:
					begin
						x1<=oldhcx-10'd80;//horizontal arm top bot
						y1<=oldhcy+9'd110;
						x2<=oldhcx-10'd80;//horizontal arm top bot
						y2<=oldhcy+9'd130;
					end
					6'd23:
					begin
						x1<=oldhcx-10'd60;//horizontal arm top bot
						y1<=oldhcy+9'd110;
						x2<=oldhcx-10'd60;
						y2<=oldhcy+9'd130;
					end
					6'd24:
					begin
						x1<=oldhcx+10'd80;//horizontal arm top
						y1<=oldhcy+9'd110;
						x2<=oldhcx+10'd60;
						y2<=oldhcy+9'd110;
					end
					6'd25:
					begin
						x1<=oldhcx+10'd80;//armleft
						y1<=oldhcy+9'd110;
						x2<=oldrcx+10'd20;
						y2<=oldrcy;
					end
					6'd26:
					begin
						x1<=oldhcx+10'd60;
						y1<=oldhcy+9'd110;
						x2<=oldrcx-10'd20;
						y2<=oldrcy;
					end
					6'd27:
					begin
						x1<=oldrcx-10'd20;
						y1<=oldrcy;
						x2<=oldrcx+10'd20;
						y2<=oldrcy;
					end
					6'd28:
					begin
						x1<=oldrcx-10'd20;
						y1<=oldrcy;
						x2<=oldrcx-10'd20;
						y2<=oldrcy-oldrcy[8:3]+10'd60;
					end
					6'd29:
					begin
						x1<=oldrcx+10'd20;
						y1<=oldrcy;
						x2<=oldrcx+10'd20;
						y2<=oldrcy-oldrcy[8:3]+10'd60;
					end
					6'd30:
					begin
						x1<=oldrcx-10'd20;
						y1<=oldrcy-oldrcy[8:3]+10'd60;
						x2<=oldrcx+10'd20;
						y2<=oldrcy-oldrcy[8:3]+10'd60;
					end
					6'd31:
					begin
						x1<=oldhcx+10'd80;//horizontal arm top bot
						y1<=oldhcy+9'd130;
						x2<=oldhcx+10'd60;
						y2<=oldhcy+9'd130;
					end
					6'd32:
					begin
						x1<=oldhcx+10'd80;//horizontal arm top bot
						y1<=oldhcy+9'd130;
						x2<=oldrcx+10'd20;
						y2<=oldrcy-oldrcy[8:3]+10'd60;					
					end
					6'd33:
					begin
						x1<=oldhcx+10'd60;
						y1<=oldhcy+9'd130;
						x2<=oldrcx-10'd20;
						y2<=oldrcy-oldrcy[8:3]+10'd60;
					end
					6'd34:
					begin
						x1<=oldhcx+10'd80;//horizontal arm top bot
						y1<=oldhcy+9'd110;
						x2<=oldhcx+10'd80;//horizontal arm top bot
						y2<=oldhcy+9'd130;
					end
					6'd35:
					begin
						x1<=oldhcx+10'd60;//horizontal arm top bot
						y1<=oldhcy+9'd110;
						x2<=oldhcx+10'd60;
						y2<=oldhcy+9'd130;
					end
					6'd36:
					begin
						x1<=oldhcx-10'd40; //body
						y1<=oldhcy+10'd110;
						x2<=oldhcx+10'd40;
						y2<=oldhcy+10'd110;
					end
					6'd37:
					begin
						x1<=oldhcx-10'd40; //body
						y1<=oldhcy+10'd110;
						x2<=oldhcx-10'd40;
						y2<=oldhcy+10'd230;
					end
					6'd38:
					begin
						x1<=oldhcx+10'd40;
						y1<=oldhcy+10'd110;
						x2<=oldhcx+10'd40;
						y2<=oldhcy+10'd230;
					end
					6'd39:
					begin
						x1<=oldhcx-10'd40;
						y1<=oldhcy+10'd230;
						x2<=oldhcx+10'd40;
						y2<=oldhcy+10'd230;
					end
					6'd40:
					begin
						x1<=oldhcx-10'd30+oldhcx[9:3]-10'd40;
						y1<=oldhcy+10'd100;
						x2<=oldhcx+10'd50+oldhcx[9:3]-10'd40;
						y2<=oldhcy+10'd100;
					end
					6'd41:
					begin
						x1<=oldhcx-10'd30+oldhcx[9:3]-10'd40;
						y1<=oldhcy+10'd100;
						x2<=oldhcx-10'd40;
						y2<=oldhcy+10'd110;
					end
					6'd42:
					begin
						x1<=oldhcx+10'd50+oldhcx[9:3]-10'd40;
						y1<=oldhcy+10'd100;
						x2<=oldhcx+10'd40;
						y2<=oldhcy+10'd110;
					end
					6'd43:
					begin
						x1<=oldhcx-10'd30+oldhcx[9:3]-10'd40;
						y1<=oldhcy+10'd100;
						x2<=oldhcx-10'd30+oldhcx[9:3]-10'd40;
						y2<=oldhcy+10'd220;
					end
					6'd44:
					begin
						x1<=oldhcx+10'd50+oldhcx[9:3]-10'd40;
						y1<=oldhcy+10'd100;
						x2<=oldhcx+10'd50+oldhcx[9:3]-10'd40;
						y2<=oldhcy+10'd220;
					end
					6'd45:
					begin
						x1<=oldhcx-10'd30+oldhcx[9:3]-10'd40;
						y1<=oldhcy+10'd220;
						x2<=oldhcx+10'd50+oldhcx[9:3]-10'd40;
						y2<=oldhcy+10'd220;
					end
					6'd46:
					begin
						x1<=oldhcx-10'd30+oldhcx[9:3]-10'd40;
						y1<=oldhcy+10'd220;
						x2<=oldhcx-10'd40;
						y2<=oldhcy+10'd230;
					end
					6'd47:
					begin
						x1<=oldhcx+10'd50+oldhcx[9:3]-10'd40;
						y1<=oldhcy+10'd220;
						x2<=oldhcx+10'd40;
						y2<=oldhcy+10'd230;
					end
				endcase
	end

endmodule
